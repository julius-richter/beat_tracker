BZh91AY&SY�BA �߀Py���g߰����`tz`f)A@s F	�0M`�L4i0S*@j4  � �R@        	)�)�?T���4y4C�mL�ڇ��z�M=A�& �4d40	�10�A&&��d*~LT�zMOMG���C�5F���(3�(���R��Pj���ѨB6 (���)���P�ʮ$D��Z%H1���:�'e{+Z�T!"��    `���#[>;�q�3��%�?�ׄ΁K�$3����I��j��KF1�#n��K���(<���BJ8Q��/]0���y��O5�&���v<���UFUw9��E_�����tӚ���Ľ�{����k>�f��R1!'��,7�a���@C��bxr����MVCb	H��H�K��+ezcb�	j���|�A�kƮ1G���,�L"je&F4�
L�V�.=�@g�m�A3#�
s��m1�ʲҭ4��b]$
��/�SU1����0��/6 �P�X�$�8ʆ\5�>W1Ne�S��2���7��j��ې��m�&��Z�{u�h�ī)���k�F��P��4�ֈ݂�&tqE��.��X�Pa�o����p�[�6�lcm�C���5��l_4P��S���ޙYɫ�NP.��%�W��l���`�*
B����-F�HGav/���&���� a��2���"�(���,�Vꔝ4�����Ҧu��x��~6)��9�U�e}):q�Q����}24Z̊0��ʽP����1
������*k�0�m�N��[!.t-f1����3|.�ZɅs�����c�[����C��B���S�O��t�X
��� 6���0h�(%�jv�	)O�VV"�ͩ^�Z��1�w���;eiR�Q���e�UȄ� ��[R��T�X�LP�J���W���}{�nk`Q"Di�Ph"V�w	��>!��hp���eY�N!d�y�p��{��ҁJ�%Ũtw�u�>g?�v�]|��M���\�CY�*�J����O�k)�u=�<�B�]a�0�?�ܐ������ z�q`�o���zC�H���x���x]������-�C�l����0�Ӛ�����8�,�,��d��jP�(��Q8!1l��E �����k����2Dh��woߐ���E=���Ap��v/IX �i<��T=�d\�%�̮�1���3)�Hp�����<�n��¤���S���)�/,��8�bsb��]�E�F�G�qQ�HLΚ��䕁�����2��o��m���=wE0�s^�a�6��RL-�u�1�<33�
u�5��a;..�mڿa�kW���̂�z=���s���NE�p/���o�'���(����b
��w$S�	
!�